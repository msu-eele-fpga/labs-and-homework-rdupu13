library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity led_pattern_generator_tb is
end entity;

architecture led_pattern_generator_tb_arch of led_pattern_generator_tb is
	
	
	
	
	begin
		
		
		
end architecture;