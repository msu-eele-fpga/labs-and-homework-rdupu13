../../hdl/pwm-rgb-led/de10nano_top.vhd