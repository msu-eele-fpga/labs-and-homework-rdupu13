../../hdl/pwm/de10nano_top.vhd