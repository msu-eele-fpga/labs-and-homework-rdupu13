library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.assert_pkg.all;
use work.print_pkg.all;
use work.tb_pkg.all;

entity async_conditioner is
	port (
		clk   : in  std_ulogic;
		rst   : in  std_ulogic;
		async : in  std_ulogic;
		sync  : out std_ulogic
	);
end entity;

architecture async_conditioner_arch of async_conditioner is
	
	
	
	begin
		
		
		
end architecture;